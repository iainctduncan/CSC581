BZh91AY&SY�lN �_�Py����߰?���P�RAT�P���A�ɓ&F�L�L0&&�	�&L�&	���`LM&L�LM2100� ��@54�=�S���  4i�ڐD�h�
z���ڞF��1� �bzC��<JQ�!���t!�pQ��)�bقI
@�\_{��T��.�K�1�xw�8Po���G�Nf�����z��1�I'&.CC���޽��TU�������c g`s����f;�ű�2�T�!��ս��%���@�i5c$
�o3b�G����ii(#��j�DoSFב��dɄ�
5�yI	�eFa0&�<�ag�zjb�`�G�l�ǁ���ذ�Ֆ43 ��j	sM='�Ӂ$(�4Q��x[lh�����<F1�I$�I$�:^�:V�9��{�d	=�=� �5������9�6A�F0���1{�	jl��� ���$$9ئP�E=���ղ���-��u?X�u��������ѫplw��C0�-����Z���|]��ƃ�Y-M�%ӡ����?�<�"��v	���"�4}P*�
��������3��K#�f�]�҇�av�h���<�C�b��Hi
��f��"=��ݤ  ��ȸf`-�d�Ǔ�I<�3���|�� ��I<�;�ƚx RH����͞!�pf���8�ڬQ�I���-HC��h��)�	W[8��j��܆a�����(X��Bq\���0��];T�C��m�u3WU5�n�����P���^����hJ5#��~���ױ�� E9��{B�h���P�S[��,o8�'�o1 u��{�0�����H�K��S�Y����u3T��눈�V�5a��B�lT�j0����,��)V�¬���,�����{F��ƈi]O<���s�[���@�=��M�C���;�|�X����&j' $��@�}^o��rn�6���̍�%��3d�c&L��� m�Ϲ��W&��4L[B��w@����c;������t���Zq�`�f#�3bb$��=K5�`�t��ShIKc�c����� ���/����9��_�]��BC	�]8