BZh91AY&SY�6�u  �_�Px����߰?���@͠ 5&�e4ѐh�4@  hz����S�0�� � h   �12dф�14�&���'��h��Bd� mOS4�a4�	���J?&��&��M���$Q�w5F���8/�:wH�ȏ�F���>�]yO͓�66�@N�}I�0�n&�N;�P��0�X�g���Z�'�«�c��:�:�k1`2z�!sj�L�<�����y�Q��"l�Օ�����9��Úɍ�sm�|{�ȹz3�R��"�﯄�N�<��Z�E�͆����d�$AXQ&p��|1��a肇�F���ԥm4�*� Ĝ����dxh�u,��D�ܚ����a0��1��� b#QY"��=�Լ�lޑ=��}3DK��A�.�/�U�&1cM�A ͫB�И]J���xIɭT$S� I��Ӟh�ĥ�eU�>\IXiMƂ{rԞ�C�e���Cx����K�0y��ҡq/��?y�Z��7*.�#��٬Ү�XW�b���o�L�b��y+�w����F���ػ���N 4ҧ�ע�1!�F#L���h8a�"��f�%3�)Zy�� k]��d��̚�SV�9Z,7�P��/��I��MiZ���Ϟ�*{q:�˰�({qӷu_�Gq��p*��l]|�A������*0D�o�J}0�jڍq����#+9n&��r���R����1�>%���$�՜?���H��]������5���F��kT��������gE����)�Y���